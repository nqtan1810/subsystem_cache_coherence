//////////////////////////////////////////////////////////////////////////////////
//
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ns

module decoder(
    input [1:0] way,
    output reg w3, w2, w1, w0
    );
    
    always @(*) begin
        case(way)
            2'b00: {w3, w2, w1, w0} = 4'b0001;
            2'b01: {w3, w2, w1, w0} = 4'b0010;
            2'b10: {w3, w2, w1, w0} = 4'b0100;
            2'b11: {w3, w2, w1, w0} = 4'b1000;
            default: {w3, w2, w1, w0} = 4'b0001;
        endcase
    end
    
endmodule
